module muxNto1 #(
    parameter N = 8,
    parameter SEL = 3     
)(
    input  [N-1:0] I,
    input  [SEL-1:0] S,
    output reg Y
);
    always @(*) begin
        Y = I[S];
    end
endmodule



/*output
meenakshi@meenakshi-Inspiron-3501:~/verilog/muxNto1$ vvp muxNto1.out
VCD info: dumpfile muxNto1.vcd opened for output.
$time=0|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=000|Y=0
$time=10|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=001|Y=0
$time=20|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=010|Y=1
$time=30|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=011|Y=1
$time=40|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=100|Y=0
$time=50|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=101|Y=1
$time=60|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=110|Y=0
$time=70|N=00000000000000000000000000001000|SEL=00000000000000000000000000000011|I=10101100|S=111|Y=1
muxNto1_tb.v:29: $finish called at 80 (1s)
*/
